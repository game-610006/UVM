class jux_axi4_virtual_sequencer extends uvm_sequencer;
`uvm_component_utils(jux_axi4_virtual_sequencer)

function new(input string name="jux_axi4_virtual_sequencer", input uvm_component parent=null);
	super.new(name, parent);
//	$display("========in virtual_seq function new=======\n");
endfunction


endclass
