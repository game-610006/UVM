`include "jux_axi4_env_pkg.sv"
import jux_axi4_env_pkg::*;

import uvm_pkg::*;
`include "jux_axi4_test.sv"
`include "test.sv"
