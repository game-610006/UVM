`ifndef JUX_DATA_WIDTH
	`define JUX_DATA_WIDTH 32
`endif

parameter int DATA_WIDTH = `JUX_DATA_WIDTH;
parameter int HM_DATA_WIDTH = `JUX_DATA_WIDTH;
